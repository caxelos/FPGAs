


`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:11:29 11/26/2016 
// Design Name: 
// Module Name:    VRAM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module greenRAM(
   input CLK,
	input SSR,//reset here
	input EN,
	input WE,
	input [13:0] ADDR_IN,
	input DATA_IN,
	output DATA_OUT
);


		
/*
 - 16Kx1 VRAM memory(single-port) 

 - I create 3 instances of that module, one for each color
 to make the 128x96MEM
*/ 

   RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("READ_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The following INIT_xx declarations specify the initial contents of the RAM
      /*
*************************   1st shape   ****************************************
      */		
		// Address 0 to 4095
		            
      .INIT_00(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//kokkino
      .INIT_01(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//aspro
      .INIT_02(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//kokkino
      .INIT_03(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//aspro
      .INIT_04(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//...
      .INIT_05(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_06(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_08(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_09(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0B(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      /*
*************************		2nd shape   ***************************************************
		*/
		.INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//prasino/aspro
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 4096 to 8191
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      /*
*************************   3rd shape   *****************************************************		
		*/
		.INIT_18(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//mple/aspro
      .INIT_19(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1A(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1B(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1C(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1E(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 8192 to 12287
      .INIT_20(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_21(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_22(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_23(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      /*
*************************   4th shape   ****************************************************
        1100_1111_1100...C_F_C_F_C_F
		  (prasino-mple-aspro-aspro-aspro-kokkino)*
		          C          F           C  
		*/		                                          
		.INIT_24(256'h00000000000000000000000000000000_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),//poluxroma
      .INIT_25(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_26(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_27(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_28(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_29(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_2A(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_2B(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_2C(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_2D(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_2E(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
      .INIT_2F(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF_00000000000000000000000000000000),
      // Address 12288 to 16383
		 /*
*************************   NO MORE MEMORY   ****************************************************
      */		
		
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),//mia mavri grammi edw
      .INIT_31(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_32(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_33(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_34(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_35(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_36(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_37(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_38(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_39(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_3A(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_3B(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_3C(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_3D(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_3E(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0),
      .INIT_3F(256'hF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0FFF0F0)
   ) RAMB16 (
      .DO(DATA_OUT),      // 1-bit Data Output
      .ADDR(ADDR_IN),  // 14-bit Address Input
      .CLK(CLK),    // Clock
      .DI(DATA_IN),      // 1-bit Data Input
      .EN(EN),      // RAM Enable Input
      .SSR(SSR),    // Synchronous Set/Reset Input
      .WE(WE)       // Write Enable Input   );
   );


endmodule
